/******************************************************************************
*
*                    Copyright 2010-2011 Dolak-NER Systems.
*                    All rights reserved worldwide.
*
*******************************************************************************/

`ifndef SDL_VERSION_DEFINES_SCH
`define SDL_VERSION_DEFINES_SCH

  `define SDL_NAME SDL
  `define SDL_MAJOR_REV 1
  `define SDL_MINOR_REV 0
  `define SDL_FIX_REV   0

  `define SDL_VERSION_STRING `"`SDL_NAME``-```SDL_MAJOR_REV``.```SDL_MINOR_REV``.```SDL_FIX_REV`"

`endif



/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/

/******************************************************************************
*
*                    Copyright 2010-2011 Dolak-NER Systems.
*                    All rights reserved worldwide.
*
*******************************************************************************/

`ifndef BASE_SVH
`define BASE_SVH
  
  `include "sdl_base/sdl_connections.svh"
  `include "sdl_base/sdl_agent_base.sv"
  `include "sdl_base/sdl_system_base.sv"
  `include "sdl_base/sdl_block_base.sv"
  `include "sdl_base/sdl_fsm_base.sv"
  `include "sdl_base/sdl_signal_base.sv"
  `include "sdl_base/sdl_process_base.sv"
  `include "sdl_base/sdl_process_input_fifo.sv"

`endif


/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/


//-----------------------------------------------------------------------------------------------
//   Copyright 2010-2011 Armen L. Khachatryan (armenkhl@gmail.com)
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//-----------------------------------------------------------------------------------------------

`ifndef PROCESS_BASE_SV
`define PROCESS_BASE_SV

`include "sdl_base/sdl_process_base.svh"


  function sdl_process_base::new(string name, uvm_component parent);
    super.new(name, parent);
    put_port = new("put_port", this);
    input_queue = new("input_queue", this);
    fsm = new("fsm", this);
  endfunction


`endif


/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/

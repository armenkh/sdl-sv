/******************************************************************************
*
*                    Copyright 2010-2011 Dolak-NER Systems.
*                    All rights reserved worldwide.
*
*******************************************************************************/

`ifndef AGENT_BASE_SV
`define AGENT_BASE_SV

class sdl_agent_base extends uvm_component;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction


endclass : sdl_agent_base

`endif


/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/

/******************************************************************************
*
*                    Copyright 2010-2011 Dolak-NER Systems.
*                    All rights reserved worldwide.
*
*******************************************************************************/

`ifndef SDL_PRINT_SVH
`define SDL_PRINT_SVH


`define sdl_info(MSG,VERBOSITY) `uvm_info("SDL-SV", MSG, VERBOSITY)

`endif

/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/

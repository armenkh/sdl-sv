//-----------------------------------------------------------------------------------------------
//   Copyright 2010-2011 Armen L. Khachatryan (armenkhl@gmail.com)
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//-----------------------------------------------------------------------------------------------

`ifndef SDL_PRINT_SVH
`define SDL_PRINT_SVH


`define sdl_info(MSG,VERBOSITY)  `uvm_info ("SDL-SV", MSG, VERBOSITY)
`define sdl_warning(MSG)         `uvm_warning ("SDL-SV", MSG)
`define sdl_error(MSG)           `uvm_error("SDL-SV", MSG)

`endif

/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/

//-----------------------------------------------------------------------------------------------
//   Copyright 2010-2011 Armen L. Khachatryan (armenkhl@gmail.com)
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//-----------------------------------------------------------------------------------------------

`ifndef SDL_VERSION_DEFINES_SCH
`define SDL_VERSION_DEFINES_SCH

  `define SDL_NAME SDL
  `define SDL_MAJOR_REV 1
  `define SDL_MINOR_REV 0
  `define SDL_FIX_REV   0

  `define SDL_VERSION_STRING `"`SDL_NAME``-```SDL_MAJOR_REV``.```SDL_MINOR_REV``.```SDL_FIX_REV`"

`endif



/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/

/******************************************************************************
*
*                    Copyright 2010-2011 Dolak-NER Systems.
*                    All rights reserved worldwide.
*
*******************************************************************************/
  

class sdl_signal_base extends uvm_transaction;

  // Function: new
  //
  // Creates a new signal object. The name is the instance name of the
  // transaction. If not supplied, then the object is unnamed.
  
  extern function new (string name="", uvm_component initiator = null);


  
endclass : sdl_signal_base


/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/



/******************************************************************************
*
*                    Copyright 2010-2011 Dolak-NER Systems.
*                    All rights reserved worldwide.
*
*******************************************************************************/

`ifndef SDL_MACROS_SVH
`define SDL_MACROS_SVH

  `include "sdl_macros/sdl_version_defines.svh"
  `include "sdl_macros/sdl_print.sv"
  
`endif


/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/

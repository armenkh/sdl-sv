/******************************************************************************
*
*                    Copyright 2010-2011 Dolak-NER Systems.
*                    All rights reserved worldwide.
*
*******************************************************************************/


  `include "sdl_pkg.svh"



/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/

/******************************************************************************
*
*                    Copyright 2010-2011 Dolak-NER Systems.
*                    All rights reserved worldwide.
*
*******************************************************************************/

`include "sdl_base/sdl_signal_base.svh"

// new
// ---


function sdl_signal_base::new (string name="", 
                               uvm_component initiator = null);
  super.new(name, initiator);
endfunction // sdl_signal_base




/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/

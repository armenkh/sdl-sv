/******************************************************************************
*
*                    Copyright 2010-2011 Dolak-NER Systems.
*                    All rights reserved worldwide.
*
*******************************************************************************/

`ifndef BLOCK_BASE_SV
`define BLOCK_BASE_SV

class sdl_block_base extends sdl_agent_base;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction


endclass : sdl_block_base

`endif



/******************************************************************************
*
* REVISION HISTORY:
*    
*******************************************************************************/
